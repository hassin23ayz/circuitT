* Title: Simulation of PV cell 
* uic = use initial condition 
.tran 0.01ms 5ms uic
.include pv.net

* Control commands
* .control
* set color0 = white ; set background as white
* set color1 = black ; set foreground as white
* run
* plot v(b)
* .endc