* Title: Half Wave Rectifier
* Analysis : Transient analysis 
.tran 1us 40ms uic
.include ex02.net

* Control commands
.control
set color0 = white ; set background as white
set color1 = black ; set foreground as white
run
plot v(a) v(b)
.endc